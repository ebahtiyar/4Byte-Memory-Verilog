library verilog;
use verilog.vl_types.all;
entity fourbytememory_vlg_vec_tst is
end fourbytememory_vlg_vec_tst;
