module andgate3(x,y,z,out);
//Three input AND gate
input x,y,z;
output out;
assign out = x & y & z;
endmodule 